//-------------------------------------------------------------------------
//      lab6_toplevel.sv                                                 --
//                                                                       --
//      Created 10-19-2017 by Po-Han Huang                               --
//                        Spring 2018 Distribution                       --
//                                                                       --
//      For use with ECE 385 Experment 6                                 --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------
module lab6_toplevel( input logic [15:0] S,
								//output logic [15:0]  PC,
                      input logic Clk, Reset, Run, Continue,
                      output logic [11:0] LED,
                      output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7,
                      output logic CE, UB, LB, OE, WE,
                      output logic [19:0] ADDR,
                      inout wire [15:0] Data);

logic [15:0] S_new;
logic Reset_o, Run_O, Continue_O;
slc3 my_slc(.*,.Reset(Reset_o), .Run(Run_O), .Continue(Continue_O), .S(S_new));
// Even though test memory is instantiated here, it will be synthesized into 
// a blank module, and will not interfere with the actual SRAM.
// Test memory is to play the role of physical SRAM in simulation.
//test_memory my_test_memory(.Reset(~Reset), .I_O(Data), .A(ADDR), .*);

sync sync_1(Clk, S, S_new);
sync sync_2(Clk, Reset, Reset_o);
sync sync_3(Clk, Run, Run_O);
sync sync_4(Clk, Continue, Continue_O);

endmodule
